`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:33:59 12/15/2020 
// Design Name: 
// Module Name:    CMP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CMP(
    input [31:0] A,
    input [31:0] B,
    output zero,
	 output isge,
	 output isgreat
    );
	 
	 assign zero = (A==B)? 1'b1 : 1'b0;
	 
	 assign isge = ($signed(A) >= $signed(0))? 1'b1 : 1'b0;
	 
	 assign isgreat = ($signed(A) > $signed(0))? 1'b1 : 1'b0;


endmodule
